module execute();
endmodule 